module partial_gen_11 (
    input logic [10:0] A,
    input logic [10:0] B,
    output logic [21:0] P0,
    output logic [21:0] P1,
    output logic [21:0] P2,
    output logic [21:0] P3,
    output logic [21:0] P4,
    output logic [21:0] P5
);

    always_comb begin
        // P0
        P0 = (!B[0] && !B[1]) ? {7'b0,1'b1,14'b0} : 
               (B[0]) ? 
                    (!B[1]) ?
                         {7'b0, !B[1], B[1], B[1], 1'b0, A} :
                         {7'b0, !B[1], B[1], B[1], 1'b1, ~A} :
                    (!B[1]) ?
                         {7'b0, !B[1], B[1], B[1], A, 1'b0}:
                         {7'b0, !B[1], B[1], B[1], ~A, 1'b1};

        // P1
        P1 = ((B[2] == B[3]) && (B[1] == B[3])) ? {6'b0, 1'b1, 1'b1, 13'b0, P0[12]} : 
               (B[2]^B[1]) ?
                    (!B[3]) ?
                         {6'b0, 1'b1, ~B[3], 1'b0, A, 1'b0, P0[12]} : 
                         {6'b0, 1'b1, ~B[3], 1'b1, ~A, 1'b0, P0[12]} : 
                    (!B[3]) ?
                         {6'b0, 1'b1, ~B[3], A, 2'b0, P0[12]}:
                         {6'b0, 1'b1, ~B[3], ~A, 1'b1, 1'b0, P0[12]};

        // P2
        P2 = ((B[4] == B[5]) && (B[3] == B[5])) ? {4'b0,1'b1, 1'b1, 13'b0, ~P1[14], 2'b0} : 
               (B[4]^B[3]) ?
                    (!B[5]) ?
                         {4'b0, 1'b1, ~B[5], 1'b0, A, 1'b0, ~P1[14], 2'b0} : 
                         {4'b0, 1'b1, ~B[5], 1'b1, ~A, 1'b0, ~P1[14], 2'b0} : 
                    (!B[5]) ?
                         {4'b0, 1'b1, ~B[5], A, 2'b0, ~P1[14], 2'b0}:
                         {4'b0, 1'b1, ~B[5], ~A, 1'b1, 1'b0, ~P1[14], 2'b0};

        // P3
        P3 = ((B[6] == B[7]) && (B[5] == B[7])) ? {2'b0, 1'b1, 1'b1, 13'b0, ~P2[16], 4'b0} : 
               (B[6]^B[5]) ?
                    (!B[7]) ?
                         {2'b0, 1'b1, ~B[7], 1'b0, A, 1'b0, ~P2[16], 4'b0} : 
                         {2'b0, 1'b1, ~B[7], 1'b1, ~A, 1'b0, ~P2[16], 4'b0} : 
                    (!B[7]) ?
                         {2'b0, 1'b1, ~B[7], A, 2'b0, ~P2[16], 4'b0}:                         
                         {2'b0, 1'b1, ~B[7], ~A, 1'b1, 1'b0, ~P2[16], 4'b0};

        // P4
        P4 = ((B[8] == B[9]) && (B[7] == B[9])) ? {1'b1, 1'b1, 13'b0, ~P3[18], 6'b0} : 
               (B[8]^B[7]) ? 
                    (!B[9]) ?
                         {1'b1, ~B[9], 1'b0, A, 1'b0, ~P3[18], 6'b0} : 
                         {1'b1, ~B[9], 1'b1, ~A, 1'b0, ~P3[18], 6'b0} : 
                    (!B[9]) ?
                         {1'b1, ~B[9], A, 2'b0, ~P3[18], 6'b0}:
                         {1'b1, ~B[9], ~A, 1'b1, 1'b0, ~P3[18], 6'b0};

        // P5
        P5 = (!B[10] && !B[9]) ? {13'b0, ~P4[20], 8'b0} : 
               (B[9] && B[10]) ? 
                    {A, 2'b0, ~P4[20], 8'b0} :
               {1'b0, A, 1'b0, ~P4[20], 8'b0};

     end
endmodule